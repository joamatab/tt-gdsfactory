VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_rc_filter
  CLASS BLOCK ;
  FOREIGN tt_rc_filter ;
  ORIGIN -1.000 -5.000 ;
  SIZE 5.000 BY 216.000 ;
END tt_rc_filter
END LIBRARY

